module Settle(

);

endmodule