module GFX(
    
);


endmodule
