module Play(

);


endmodule