module Chess(

);





endmodule