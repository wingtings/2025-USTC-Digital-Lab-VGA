module Menu(
    
);





endmodule