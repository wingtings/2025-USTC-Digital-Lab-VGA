module Selector(

);

endmodule