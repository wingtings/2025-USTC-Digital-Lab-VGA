// 游戏结束逻辑判断模块, 接收 board_data, 输出 game_over 信号
module Over(
    input clkk,
    input rstn,
    input board_data [12*64-1:0],
    output reg [1:0] game_over
);







endmodule